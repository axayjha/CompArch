module notgate(A,B);
	input A;
	output B;
	assign A=!B;
endmodule
